netcdf gwf_chd01 {
dimensions:
	LINELENGTH = 300 ;
	LENAUXNAME = 16 ;
	LENBOUNDNAME = 40 ;
	NPER = 1 ;
	NLAY = 1 ;
	NROW = 1 ;
	NCOL = 100 ;
	NCPL = 100 ;
	NCELLDIM = 3 ;
	dim_chd-1_maxbound = 2 ;
	dim_chd-1_niper = 1 ;
variables:
	int dis_nlay ;
		dis_nlay:mf6_input = "DIS6:GWF_CHD01/DIS/NLAY" ;
	int dis_nrow ;
		dis_nrow:mf6_input = "DIS6:GWF_CHD01/DIS/NROW" ;
	int dis_ncol ;
		dis_ncol:mf6_input = "DIS6:GWF_CHD01/DIS/NCOL" ;
	double dis_delr(NCOL) ;
		dis_delr:_FillValue = 3.e+30 ;
		dis_delr:mf6_input = "DIS6:GWF_CHD01/DIS/DELR" ;
	double dis_delc(NROW) ;
		dis_delc:_FillValue = 3.e+30 ;
		dis_delc:mf6_input = "DIS6:GWF_CHD01/DIS/DELC" ;
	double dis_top(NLAY, NROW, NCOL) ;
		dis_top:_FillValue = 3.e+30 ;
		dis_top:mf6_input = "DIS6:GWF_CHD01/DIS/TOP" ;
	double dis_botm(NLAY, NROW, NCOL) ;
		dis_botm:_FillValue = 3.e+30 ;
		dis_botm:mf6_input = "DIS6:GWF_CHD01/DIS/BOTM" ;
	int dis_idomain(NLAY, NROW, NCOL) ;
		dis_idomain:_FillValue = -2147483647 ;
		dis_idomain:mf6_input = "DIS6:GWF_CHD01/DIS/IDOMAIN" ;
	double ic_strt(NLAY, NROW, NCOL) ;
		ic_strt:_FillValue = 3.e+30 ;
		ic_strt:mf6_input = "IC6:GWF_CHD01/IC/STRT" ;
	int npf_save_specific_discharge ;
		npf_save_specific_discharge:mf6_input = "NPF6:GWF_CHD01/NPF/SAVE_SPECIFIC_DISCHARGE" ;
	int npf_icelltype(NLAY, NROW, NCOL) ;
		npf_icelltype:_FillValue = -2147483647 ;
		npf_icelltype:mf6_input = "NPF6:GWF_CHD01/NPF/ICELLTYPE" ;
	double npf_k(NLAY, NROW, NCOL) ;
		npf_k:_FillValue = 3.e+30 ;
		npf_k:mf6_input = "NPF6:GWF_CHD01/NPF/K" ;
	double npf_k33(NLAY, NROW, NCOL) ;
		npf_k33:_FillValue = 3.e+30 ;
		npf_k33:mf6_input = "NPF6:GWF_CHD01/NPF/K33" ;
	int chd-1_print_flows ;
		chd-1_print_flows:mf6_input = "CHD6:GWF_CHD01/CHD-1/PRINT_FLOWS" ;
	int chd-1_maxbound ;
		chd-1_maxbound:mf6_input = "CHD6:GWF_CHD01/CHD-1/MAXBOUND" ;
	int chd-1_cellid(dim_chd-1_niper, dim_chd-1_maxbound, NCELLDIM) ;
		chd-1_cellid:_FillValue = -2147483647 ;
		chd-1_cellid:mf6_input = "CHD6:GWF_CHD01/CHD-1/CELLID" ;
	double chd-1_head(dim_chd-1_niper, dim_chd-1_maxbound) ;
		chd-1_head:_FillValue = 3.e+30 ;
		chd-1_head:mf6_input = "CHD6:GWF_CHD01/CHD-1/HEAD" ;
	int chd-1_iper(dim_chd-1_niper) ;
		chd-1_iper:_FillValue = -2147483647 ;
		chd-1_iper:mf6_input = "CHD6:GWF_CHD01/CHD-1/IPER" ;

// global attributes:
		:description = "MODFLOW 6 NetCDF4 file prototype" ;
		:history = "Created Thu Feb 29 15:52:48 2024" ;
		:source = "flopy v3.5.0.dev0" ;
		:mf6_modeltype = "GWF6" ;
		:mf6_modelname = "GWF_CHD01" ;
		:Conventions = "" ;
data:

 dis_nlay = 1 ;

 dis_nrow = 1 ;

 dis_ncol = 100 ;

 dis_delr = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1 ;

 dis_delc = 1 ;

 dis_top =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 dis_botm =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 dis_idomain =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 ic_strt =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 npf_save_specific_discharge = 1 ;

 npf_icelltype =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 npf_k =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 npf_k33 =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 chd-1_print_flows = 1 ;

 chd-1_maxbound = 2 ;

 chd-1_cellid =
  1, 1, 1,
  1, 1, 100 ;

 chd-1_head =
  1, 0 ;

 chd-1_iper = 1 ;
}
